`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: USTC ESLAB
// Engineer: Huang Yifan (hyf15@mail.ustc.edu.cn)
// 
// Design Name: RV32I Core
// Module Name: Write-back Data seg reg
// Tool Versions: Vivado 2017.4.1
// Description: Write-back data seg reg for MEM\WB
// 
//////////////////////////////////////////////////////////////////////////////////


//  ???��??��?????
    // MEM\WB?????????????????��??��???
    // ????????��????????????Data Extension?��?Data Cache��???????��?��????
// ��?��?��?
    // clk               ?��?����??????��
    // wb_select         �����?????????????????��?????��???????????????0?????????ALU��????��??��???????????????1?????????Memory��????�C?????��???
    // load_type         load?????��?��????
    // write_en          Data Cache??????��??
    // debug_write_en    Data Cache debug??????��??
    // addr              Data Cache????????��??��?????????ALU???��????��??��???
    // debug_addr        Data Cache???debug?????��???
    // in_data           Data Cache???????��???��???
    // debug_in_data     Data Cache???debug????��???��???
    // bubbleW           WB��????????bubble?????��
    // flushW            WB��????????flush?????��
// ��?��???
    // debug_out_data    Data Cache???debug��???????��???
    // data_WB           ?? ????????��????��?????????????????????��??��???
// ???��??��???��?  
    // ?�� ��?��????��?

module WB_Data_WB(
    input wire clk, rst, bubbleW, flushW,
    input wire wb_select,
    input wire [2:0] load_type,
    input  [3:0] write_en, debug_write_en,
    input  [31:0] addr,
    input  [31:0] debug_addr,
    input  [31:0] in_data, debug_in_data,
    output wire [31:0] debug_out_data,
    output wire [31:0] data_WB,
    output miss, ref_signal
    );

    wire [31:0] data_raw;
    wire [31:0] data_WB_raw;
    wire n_write_en;
    assign n_write_en = (write_en == 4'b1111) ? 1'b1 : 1'b0;


    /* DataCache DataCache1(
        .clk(clk),
        .write_en(write_en << addr[1:0]),
        .debug_write_en(debug_write_en),
        .addr(addr[31:2]),
        .debug_addr(debug_addr[31:2]),
        .in_data(in_data << (8 * addr[1:0])),
        .debug_in_data(debug_in_data),
        .out_data(data_raw),
        .debug_out_data(debug_out_data)
    ); */
    cache cache1 (
        .clk(clk),
        .rst(rst),
        .addr(addr),
        .wr_data(in_data),
        .rd_req(wb_select),
        .wr_req(n_write_en),
        .rd_data(data_raw),
        .miss(miss),
        .ref_signal(ref_signal)
    );
    // Add flush and bubble support
    // if chip not enabled, output output last read result
    // else if chip clear, output 0
    // else output values from cache

    reg bubble_ff = 1'b0;
    reg flush_ff = 1'b0;
    reg wb_select_old = 0;
    reg [31:0] data_WB_old = 32'b0;
    reg [31:0] addr_old;
    reg [2:0] load_type_old;

    DataExtend DataExtend1(
        .data(data_raw),
        .addr(addr_old[1:0]),
        .load_type(load_type_old),
        .dealt_data(data_WB_raw)
    );

    always@(posedge clk)
    begin
        bubble_ff <= bubbleW;
        flush_ff <= flushW;
        data_WB_old <= data_WB;
        addr_old <= addr;
        wb_select_old <= wb_select;
        load_type_old <= load_type;
    end

    assign data_WB = bubble_ff ? data_WB_old :
                                 (flush_ff ? 32'b0 : 
                                             (wb_select_old ? data_WB_raw :
                                                          addr_old));






    
endmodule